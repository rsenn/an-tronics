Amplifier
C1 9 2 100µF IC=0
D2 4 6 DI_1N4001
D1 5 4 DI_1N4001
R3 5 2 330
R2 1 2 100
C2 0 1 220µF IC=0
R4 1 10 22
C3 3 7 1µF IC=0

*SRC=1N4001;DI_1N4001;Diodes;Si;  50.0V  1.00A  3.00us   Diodes, Inc. diode
.MODEL DI_1N4001 D  ( IS=76.9p RS=42.0m BV=50.0 IBV=5.00u CJO=39.8p  M=0.333 N=1.45 TT=4.32u )

.TRAN 1ms 100ms
* .AC DEC 100 100 1MEG
.END
